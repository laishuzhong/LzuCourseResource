`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2021/09/17 16:14:49
// Design Name: 
// Module Name: float_adder_addition
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


//top file
module Floating_Point_Addition(clk,reset,x,y, result);
input clk,reset;
input [31:0] x,y;    
output [31:0] result;
//???????????????
wire[8:0] exp_diff; //????????????
wire mux_1_en; //???1 ????
wire mux_2_en; //???2 ????
wire mux_3_en; //???3 ????
wire[7:0] mux_1_output; //???1 ?????
wire[31:0] mux_2_output; //???2 ?????
wire[31:0] mux_3_output; //???3 ?????
wire[7:0] shift_right_bit; //????????????????
wire[26:0] shift_right_output; //?????????

wire[27:0] big_alu_result; //????????????
wire[7:0] shift_right_bits; //?????????????
wire[7:0] shift_left_bits; //?????????????
wire shift_right_en; //???????????????
wire shift_left_en; //???????????????
wire[27:0] mux_4_output; //???4 ?????
wire mux_4_en; //???4 ????
wire[27:0] shift_left_right_output; //??????????????????
wire[7:0] incre_bit; //??????????
wire[7:0] decre_bit; //??????????
wire incre_en; //????????????
wire decre_en; //????????????
wire mux_5_en; //???5 ????
wire[7:0] mux_5_output; //???5 ?????
wire[7:0] rounding_exp_result; //????????????
wire[8:0] incre_decre_output; //??????????????
wire[27:0] fra_result; //????
//wire[31:0] result;
wire overflow; //?????

//?????????????????
Small_Alu
Small_Alu_instance(
//????
clk,
reset,
x,
y,
//????
exp_diff //????????????????
);

//???
Control
Control_instance(
clk,
reset,
exp_diff,
big_alu_result,
fra_result,
shift_right_bits,

shift_left_bits,
shift_right_en,
shift_left_en,
shift_right_bit,
incre_bit,
decre_bit,
incre_en,
decre_en,
mux_1_en,
mux_2_en,
mux_3_en,
mux_4_en,
mux_5_en
);

//???1
Mux_1
Mux_1_instance(
clk,
reset,
x,
y,
mux_1_en,
mux_1_output
);

//???2
Mux_2
Mux_2_instance(
clk,
reset,
x,
y,
mux_2_en,
mux_2_output
);

//???3
Mux_3
Mux_3_instance(
clk,
reset,
x,
y,
mux_3_en,
mux_3_output
);

Shift_Right //????????????????
Shift_Right_instance(
clk,
reset,
shift_right_bit,
mux_2_output,
shift_right_output //??shift_right_bit??mux_2_output ????
);

//???????????
Big_Alu
Big_Alu_instance(
clk,
reset,
shift_right_output,
mux_3_output,
big_alu_result //mux_3_output ?shift_right_output ????????big_alu_result
);

//???4
Mux_4
Mux_4_instance(
clk,
reset,
mux_4_en,
big_alu_result,
fra_result,
mux_4_output
);

Shift_Left_Right //???????????
Shift_Left_Right_instance(
clk,
reset,
shift_left_bits,
shift_right_bits,
shift_left_en,
shift_right_en,
mux_4_output,
shift_left_right_output
);

//???5
Mux_5
Mux_5_instance(
clk,
reset,
mux_5_en,
mux_1_output,
rounding_exp_result,
mux_5_output
);

Incre_Decre //???????????
Incre_Decre_instance(
clk,
reset,
incre_bit,
decre_bit,
incre_en,
decre_en,
mux_5_output,
incre_decre_output //??incre_bit ?incre_en??mux_5_output??????decre_bit ?decre_en??mux_5_output ???
);

//??????
Rounding
Rounding_instance(
clk,
reset,
shift_left_right_output,
incre_decre_output,
rounding_exp_result,
fra_result, //????
result,
overflow //????
);

endmodule
